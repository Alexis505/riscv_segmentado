module imem(input logic  [31:0] a,
	    output logic [31:0] rd);

	logic [31:0] RAM[63:0]; //arreglo de 64 filas de 32 bits cada una
	
	initial 
		$readmemh("riscvtest.txt",RAM);

	assign rd = RAM[a[31:2]]; //word aligned

endmodule



//	*************************
//      * 			*
//  --->* A			*
//	*			*
//	*	Instruction	*
//	*	Memory		*
//	*			*
//	*			*
//	*			*
//  <---* RD			*
//	*			*
//	*************************
